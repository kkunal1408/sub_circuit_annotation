MACRO CMC_NMOS_S_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_S_n12_X3_Y1 0 0 ;
  SIZE 3.8400 BY 1.5120 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.6600 0.0480 1.7000 0.4560 ;
      LAYER M3 ;
        RECT 1.9800 0.0480 2.0200 0.4560 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.7400 0.1320 1.7800 0.5400 ;
      LAYER M3 ;
        RECT 2.0600 0.1320 2.1000 0.5400 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.8200 0.2160 1.8600 0.6240 ;
      LAYER M3 ;
        RECT 2.1400 0.2160 2.1800 0.6240 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.9000 0.3000 1.9400 0.7080 ;
      LAYER M3 ;
        RECT 2.2200 0.3000 2.2600 0.7080 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 3.8040 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 1.0560 0.9760 1.2960 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 1.0560 1.6160 1.2960 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 1.0560 2.2560 1.2960 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 1.0560 2.8960 1.2960 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 1.0560 3.5360 1.2960 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 3.4760 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.4040 3.4760 0.4360 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 2.9960 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.4880 2.9960 0.5200 ;
    LAYER M2 ;
      RECT 1.0040 0.2360 3.6360 0.2680 ;
    LAYER M2 ;
      RECT 1.0040 0.5720 3.6360 0.6040 ;
    LAYER M2 ;
      RECT 0.2840 0.3200 3.5560 0.3520 ;
    LAYER M2 ;
      RECT 0.2840 0.6560 3.5560 0.6880 ;
  END
END CMC_NMOS_S_n12_X3_Y1
MACRO CMC_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN CMC_NMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 1.5120 ;
  PIN SA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 2.3560 0.1000 ;
    END
  END SA
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.1960 0.1840 ;
    END
  END DA
  PIN SB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.8440 0.2360 1.7160 0.2680 ;
    END
  END SB
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.3200 1.5560 0.3520 ;
    END
  END DB
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.4040 2.2760 0.4360 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 2.5240 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 1.0560 0.9760 1.2960 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 1.0560 1.6160 1.2960 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 1.0560 2.2560 1.2960 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
  END
END CMC_NMOS_n12_X2_Y1
MACRO DCL_NMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 1.5120 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.0480 0.2600 0.2880 ;
      LAYER M3 ;
        RECT 0.3800 0.0480 0.4200 0.2880 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.1320 0.3400 0.3720 ;
      LAYER M3 ;
        RECT 0.4600 0.1320 0.5000 0.3720 ;
    END
  END D
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 0.6040 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.2360 0.4360 0.2680 ;
    LAYER M2 ;
      RECT 0.2040 0.1520 0.5160 0.1840 ;
    LAYER M2 ;
      RECT 0.2040 0.3200 0.5160 0.3520 ;
  END
END DCL_NMOS_n12_X1_Y1
MACRO DCL_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 1.5120 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.5400 0.0480 0.5800 0.2880 ;
      LAYER M3 ;
        RECT 0.7000 0.0480 0.7400 0.2880 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.1320 0.6600 0.3720 ;
      LAYER M3 ;
        RECT 0.7800 0.1320 0.8200 0.3720 ;
    END
  END D
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 1.2440 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 1.0560 0.9760 1.2960 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.2360 0.9160 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 1.0760 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.3200 1.0760 0.3520 ;
  END
END DCL_NMOS_n12_X2_Y1
MACRO DCL_PMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN DCL_PMOS_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 1.5120 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.0480 0.2600 0.2880 ;
      LAYER M3 ;
        RECT 0.3800 0.0480 0.4200 0.2880 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.1320 0.3400 0.3720 ;
      LAYER M3 ;
        RECT 0.4600 0.1320 0.5000 0.3720 ;
    END
  END D
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 0.6040 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.2360 0.4360 0.2680 ;
    LAYER M2 ;
      RECT 0.2040 0.1520 0.5160 0.1840 ;
    LAYER M2 ;
      RECT 0.2040 0.3200 0.5160 0.3520 ;
  END
END DCL_PMOS_n12_X1_Y1
MACRO DP_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_n12_X3_Y1 0 0 ;
  SIZE 3.8400 BY 1.5120 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2040 0.0680 3.4760 0.1000 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3640 0.1520 2.9960 0.1840 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.0040 0.2360 3.6360 0.2680 ;
    END
  END DB
  PIN GA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.2840 0.3200 2.9160 0.3520 ;
    END
  END GA
  PIN GB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.9240 0.4040 3.5560 0.4360 ;
    END
  END GB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 3.8040 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 1.0560 0.9760 1.2960 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 1.0560 1.6160 1.2960 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 1.0560 2.2560 1.2960 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 1.0560 2.8960 1.2960 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 0.0480 3.5360 0.7080 ;
    LAYER M1 ;
      RECT 3.5040 1.0560 3.5360 1.2960 ;
    LAYER M1 ;
      RECT 3.4240 0.0480 3.4560 0.7080 ;
    LAYER M1 ;
      RECT 3.5840 0.0480 3.6160 0.7080 ;
  END
END DP_NMOS_n12_X3_Y1
MACRO SCM_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_n12_X2_Y1 0 0 ;
  SIZE 2.5600 BY 1.5120 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.1000 0.0480 1.1400 0.3720 ;
      LAYER M3 ;
        RECT 1.3400 0.0480 1.3800 0.3720 ;
    END
  END S
  PIN DA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.1800 0.1320 1.2200 0.4560 ;
      LAYER M3 ;
        RECT 1.4200 0.1320 1.4600 0.4560 ;
    END
  END DA
  PIN DB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.2600 0.2160 1.3000 0.5400 ;
      LAYER M3 ;
        RECT 1.5000 0.2160 1.5400 0.5400 ;
    END
  END DB
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 2.5240 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 1.0560 0.9760 1.2960 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 1.0560 1.6160 1.2960 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 1.0560 2.2560 1.2960 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 2.3560 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.3200 2.3560 0.3520 ;
    LAYER M2 ;
      RECT 0.2840 0.1520 2.2760 0.1840 ;
    LAYER M2 ;
      RECT 0.2840 0.4040 2.2760 0.4360 ;
    LAYER M2 ;
      RECT 1.0040 0.2360 1.5560 0.2680 ;
    LAYER M2 ;
      RECT 1.0040 0.4880 1.5560 0.5200 ;
  END
END SCM_NMOS_n12_X2_Y1
MACRO Switch_NMOS_n12_X2_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X2_Y1 0 0 ;
  SIZE 1.2800 BY 1.5120 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4600 0.0480 0.5000 0.3720 ;
      LAYER M3 ;
        RECT 0.7000 0.0480 0.7400 0.3720 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.5400 0.1320 0.5800 0.4560 ;
      LAYER M3 ;
        RECT 0.7800 0.1320 0.8200 0.4560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.6200 0.2160 0.6600 0.5400 ;
      LAYER M3 ;
        RECT 0.8600 0.2160 0.9000 0.5400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 1.2440 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 1.0560 0.9760 1.2960 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 0.9160 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.3200 0.9160 0.3520 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.0760 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.4040 1.0760 0.4360 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 0.9960 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.4880 0.9960 0.5200 ;
  END
END Switch_NMOS_n12_X2_Y1
MACRO Switch_NMOS_n12_X3_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_n12_X3_Y1 0 0 ;
  SIZE 1.9200 BY 1.5120 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.7800 0.0480 0.8200 0.3720 ;
      LAYER M3 ;
        RECT 1.0200 0.0480 1.0600 0.3720 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.8600 0.1320 0.9000 0.4560 ;
      LAYER M3 ;
        RECT 1.1000 0.1320 1.1400 0.4560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.9400 0.2160 0.9800 0.5400 ;
      LAYER M3 ;
        RECT 1.1800 0.2160 1.2200 0.5400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 1.8840 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 1.0560 0.9760 1.2960 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 1.0560 1.6160 1.2960 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 1.5560 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.3200 1.5560 0.3520 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 1.7160 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.4040 1.7160 0.4360 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 1.6360 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.4880 1.6360 0.5200 ;
  END
END Switch_NMOS_n12_X3_Y1
MACRO Switch_PMOS_n12_X1_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X1_Y1 0 0 ;
  SIZE 0.6400 BY 1.5120 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.1400 0.0480 0.1800 0.3720 ;
      LAYER M3 ;
        RECT 0.3800 0.0480 0.4200 0.3720 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.2200 0.1320 0.2600 0.4560 ;
      LAYER M3 ;
        RECT 0.4600 0.1320 0.5000 0.4560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.3000 0.2160 0.3400 0.5400 ;
      LAYER M3 ;
        RECT 0.5400 0.2160 0.5800 0.5400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 0.6040 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M2 ;
      RECT 0.1240 0.0680 0.4360 0.1000 ;
    LAYER M2 ;
      RECT 0.1240 0.3200 0.4360 0.3520 ;
    LAYER M2 ;
      RECT 0.2040 0.1520 0.5160 0.1840 ;
    LAYER M2 ;
      RECT 0.2040 0.4040 0.5160 0.4360 ;
    LAYER M2 ;
      RECT 0.2040 0.2360 0.5960 0.2680 ;
    LAYER M2 ;
      RECT 0.2040 0.4880 0.5960 0.5200 ;
  END
END Switch_PMOS_n12_X1_Y1
MACRO Switch_PMOS_n12_X5_Y1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X5_Y1 0 0 ;
  SIZE 3.2000 BY 1.5120 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.4200 0.0480 1.4600 0.3720 ;
      LAYER M3 ;
        RECT 1.6600 0.0480 1.7000 0.3720 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.5000 0.1320 1.5400 0.4560 ;
      LAYER M3 ;
        RECT 1.7400 0.1320 1.7800 0.4560 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.5800 0.2160 1.6200 0.5400 ;
      LAYER M3 ;
        RECT 1.8200 0.2160 1.8600 0.5400 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 1.1600 3.1640 1.1920 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 1.0560 0.3360 1.2960 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 1.0560 0.9760 1.2960 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 1.0560 1.6160 1.2960 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 1.0560 2.2560 1.2960 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 1.0560 2.8960 1.2960 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 2.8360 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.3200 2.8360 0.3520 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 2.9960 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.4040 2.9960 0.4360 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 2.9160 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.4880 2.9160 0.5200 ;
  END
END Switch_PMOS_n12_X5_Y1
MACRO Switch_PMOS_n12_X5_Y2
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_n12_X5_Y2 0 0 ;
  SIZE 3.2000 BY 2.3520 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.4200 0.0480 1.4600 1.2120 ;
      LAYER M3 ;
        RECT 1.6600 0.0480 1.7000 1.2120 ;
    END
  END S
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.5000 0.1320 1.5400 1.2960 ;
      LAYER M3 ;
        RECT 1.7400 0.1320 1.7800 1.2960 ;
    END
  END D
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.5800 0.2160 1.6200 1.3800 ;
      LAYER M3 ;
        RECT 1.8200 0.2160 1.8600 1.3800 ;
    END
  END G
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0360 2.0000 3.1640 2.0320 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.3040 0.0480 0.3360 0.7080 ;
    LAYER M1 ;
      RECT 0.3040 0.8880 0.3360 1.5480 ;
    LAYER M1 ;
      RECT 0.3040 1.8960 0.3360 2.1360 ;
    LAYER M1 ;
      RECT 0.2240 0.0480 0.2560 0.7080 ;
    LAYER M1 ;
      RECT 0.2240 0.8880 0.2560 1.5480 ;
    LAYER M1 ;
      RECT 0.3840 0.0480 0.4160 0.7080 ;
    LAYER M1 ;
      RECT 0.3840 0.8880 0.4160 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 0.0480 0.9760 0.7080 ;
    LAYER M1 ;
      RECT 0.9440 0.8880 0.9760 1.5480 ;
    LAYER M1 ;
      RECT 0.9440 1.8960 0.9760 2.1360 ;
    LAYER M1 ;
      RECT 0.8640 0.0480 0.8960 0.7080 ;
    LAYER M1 ;
      RECT 0.8640 0.8880 0.8960 1.5480 ;
    LAYER M1 ;
      RECT 1.0240 0.0480 1.0560 0.7080 ;
    LAYER M1 ;
      RECT 1.0240 0.8880 1.0560 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 0.0480 1.6160 0.7080 ;
    LAYER M1 ;
      RECT 1.5840 0.8880 1.6160 1.5480 ;
    LAYER M1 ;
      RECT 1.5840 1.8960 1.6160 2.1360 ;
    LAYER M1 ;
      RECT 1.5040 0.0480 1.5360 0.7080 ;
    LAYER M1 ;
      RECT 1.5040 0.8880 1.5360 1.5480 ;
    LAYER M1 ;
      RECT 1.6640 0.0480 1.6960 0.7080 ;
    LAYER M1 ;
      RECT 1.6640 0.8880 1.6960 1.5480 ;
    LAYER M1 ;
      RECT 2.2240 0.0480 2.2560 0.7080 ;
    LAYER M1 ;
      RECT 2.2240 0.8880 2.2560 1.5480 ;
    LAYER M1 ;
      RECT 2.2240 1.8960 2.2560 2.1360 ;
    LAYER M1 ;
      RECT 2.1440 0.0480 2.1760 0.7080 ;
    LAYER M1 ;
      RECT 2.1440 0.8880 2.1760 1.5480 ;
    LAYER M1 ;
      RECT 2.3040 0.0480 2.3360 0.7080 ;
    LAYER M1 ;
      RECT 2.3040 0.8880 2.3360 1.5480 ;
    LAYER M1 ;
      RECT 2.8640 0.0480 2.8960 0.7080 ;
    LAYER M1 ;
      RECT 2.8640 0.8880 2.8960 1.5480 ;
    LAYER M1 ;
      RECT 2.8640 1.8960 2.8960 2.1360 ;
    LAYER M1 ;
      RECT 2.7840 0.0480 2.8160 0.7080 ;
    LAYER M1 ;
      RECT 2.7840 0.8880 2.8160 1.5480 ;
    LAYER M1 ;
      RECT 2.9440 0.0480 2.9760 0.7080 ;
    LAYER M1 ;
      RECT 2.9440 0.8880 2.9760 1.5480 ;
    LAYER M2 ;
      RECT 0.2040 0.0680 2.8360 0.1000 ;
    LAYER M2 ;
      RECT 0.2040 0.3200 2.8360 0.3520 ;
    LAYER M2 ;
      RECT 0.3640 0.1520 2.9960 0.1840 ;
    LAYER M2 ;
      RECT 0.3640 0.4040 2.9960 0.4360 ;
    LAYER M2 ;
      RECT 0.2840 0.2360 2.9160 0.2680 ;
    LAYER M2 ;
      RECT 0.2840 0.4880 2.9160 0.5200 ;
    LAYER M2 ;
      RECT 0.2040 0.9080 2.8360 0.9400 ;
    LAYER M2 ;
      RECT 0.2040 1.1600 2.8360 1.1920 ;
    LAYER M2 ;
      RECT 0.3640 0.9920 2.9960 1.0240 ;
    LAYER M2 ;
      RECT 0.3640 1.2440 2.9960 1.2760 ;
    LAYER M2 ;
      RECT 0.2840 1.0760 2.9160 1.1080 ;
    LAYER M2 ;
      RECT 0.2840 1.3280 2.9160 1.3600 ;
  END
END Switch_PMOS_n12_X5_Y2
